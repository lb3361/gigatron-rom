sd-default.vhd